//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.12
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Fri Oct 24 19:53:59 2025

module font8x8 (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [10:0] ad;

wire [23:0] prom_inst_0_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[23:0],dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 8;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h006C6CFE6CFE6C6C0000000000006C6C00180018183C3C180000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000C060600076CCDC76386C3800C6663018CCC6000030F80C78C07C30;
defparam prom_inst_0.INIT_RAM_0A = 256'h00003030FC3030000000663CFF3C660000603018181830600018306060603018;
defparam prom_inst_0.INIT_RAM_0B = 256'h0080C06030180C06003030000000000000000000FC0000006030300000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0078CC0C380CCC7800FCCC60380CCC7800FC303030307030007CE6F6DECEC67C;
defparam prom_inst_0.INIT_RAM_0D = 256'h00303030180CCCFC0078CCCCF8C060380078CC0C0CF8C0FC001E0CFECC6C3C1C;
defparam prom_inst_0.INIT_RAM_0E = 256'h603030000030300000303000003030000070180C7CCCCC780078CCCC78CCCC78;
defparam prom_inst_0.INIT_RAM_0F = 256'h00300030180CCC78006030180C1830600000FC0000FC000000183060C0603018;
defparam prom_inst_0.INIT_RAM_10 = 256'h003C66C0C0C0663C00FC66667C6666FC00CCCCFCCCCC78300078C0DEDEDEC67C;
defparam prom_inst_0.INIT_RAM_11 = 256'h003E66CEC0C0663C00F06068786862FE00FE6268786862FE00F86C6666666CF8;
defparam prom_inst_0.INIT_RAM_12 = 256'h00E6666C786C66E60078CCCC0C0C0C1E007830303030307800CCCCCCFCCCCCCC;
defparam prom_inst_0.INIT_RAM_13 = 256'h00386CC6C6C66C3800C6C6CEDEF6E6C600C6C6D6FEFEEEC600FE6662606060F0;
defparam prom_inst_0.INIT_RAM_14 = 256'h0078CC1C70E0CC7800E6666C7C6666FC001C78DCCCCCCC7800F060607C6666FC;
defparam prom_inst_0.INIT_RAM_15 = 256'h00C6EEFED6C6C6C6003078CCCCCCCCCC00FCCCCCCCCCCCCC007830303030B4FC;
defparam prom_inst_0.INIT_RAM_16 = 256'h007860606060607800FE6632188CC6FE0078303078CCCCCC00C66C38386CC6C6;
defparam prom_inst_0.INIT_RAM_17 = 256'hFF0000000000000000000000C66C381000781818181818780002060C183060C0;
defparam prom_inst_0.INIT_RAM_18 = 256'h0078CCC0CC78000000DC66667C6060E00076CC7C0C7800000000000000183030;
defparam prom_inst_0.INIT_RAM_19 = 256'hF80C7CCCCC76000000F06060F0606C380078C0FCCC7800000076CCCC7C0C0C1C;
defparam prom_inst_0.INIT_RAM_1A = 256'h00E66C786C6660E078CCCC0C0C0C000C007830303070003000E66666766C60E0;
defparam prom_inst_0.INIT_RAM_1B = 256'h0078CCCCCC78000000CCCCCCCCF8000000C6D6FEFECC00000078303030303070;
defparam prom_inst_0.INIT_RAM_1C = 256'h00F80C78C07C000000F0606676DC00001E0C7CCCCC760000F0607C6666DC0000;
defparam prom_inst_0.INIT_RAM_1D = 256'h006CFEFED6C60000003078CCCCCC00000076CCCCCCCC000000183430307C3010;
defparam prom_inst_0.INIT_RAM_1E = 256'h001C3030E030301C00FC643098FC0000F80C7CCCCCCC000000C66C386CC60000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000DC7600E030301C3030E00018181800181818;
defparam prom_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_28 = 256'h00FCE660F0646C3818187EC0C07E181800181818180018180000000000000000;
defparam prom_inst_0.INIT_RAM_29 = 256'h78CC386C6C38633E00181818001818183030FC30FC78CCCC00C67C6C7CC60000;
defparam prom_inst_0.INIT_RAM_2A = 256'h00003366CC663300000000003E6C6C3C3C4299A1A199423C00000000000000CC;
defparam prom_inst_0.INIT_RAM_2B = 256'h000000000000007E3C42A5B9A5B9423C000000000000000000000C0CFC000000;
defparam prom_inst_0.INIT_RAM_2C = 256'h000000380C180C380000003C30180C38007E0018187E181800000000386C6C38;
defparam prom_inst_0.INIT_RAM_2D = 256'h0000001818000000001B1B1B7BDBDB7FC0607C66666600000000000000003018;
defparam prom_inst_0.INIT_RAM_2E = 256'h0000CC663366CC0000000000386C6C380000000038103010780C180000000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h0078CCC060300030016735DB2DC623C00FCC6633DECCC6C3C0CF6F37BDCCC6C3;
defparam prom_inst_0.INIT_RAM_30 = 256'h00C6FEC67C00DC7600C6FEC67C006C3800C6FEC66C38000E00C6FEC66C3800E0;
defparam prom_inst_0.INIT_RAM_31 = 256'h780C1878CCC0CC7800CECCCCFECC6C3E00CCFCCC7800303000C6C6FEC66C38C6;
defparam prom_inst_0.INIT_RAM_32 = 256'h00FC607860FC006C00FC607860FC483000FC607860FC001C00FC607860FC00E0;
defparam prom_inst_0.INIT_RAM_33 = 256'h00783030307800CC0078303078004830007830303078001C00783030307800E0;
defparam prom_inst_0.INIT_RAM_34 = 256'h00183C663C18000E00183C663C18007000CCDCFCECCC00FC00FC6666F6F666FC;
defparam prom_inst_0.INIT_RAM_35 = 256'h00006C3810386C0000183C66663C18C3007CC6C67C00DC7600183C663C18663C;
defparam prom_inst_0.INIT_RAM_36 = 256'h003C66666600663C003C66666666000E003C66666666007000B86CF6DECE6C3A;
defparam prom_inst_0.INIT_RAM_37 = 256'hC0C0F8CCF8CC7800F0607C66667C60F00018183C6666000E0078CCCCCCCC00CC;
defparam prom_inst_0.INIT_RAM_38 = 256'h007ECC7C0C78DC76003F663E063CC37E007ECC7C0C78001C007ECC7C0C7800E0;
defparam prom_inst_0.INIT_RAM_39 = 256'h380C78C0C0780000007FCC7F0C7F0000007ECC7C0C783030007ECC7C0C7800CC;
defparam prom_inst_0.INIT_RAM_3A = 256'h0078C0FCCC7800CC003C607E663CC37E0078C0FCCC78001C0078C0FCCC7800E0;
defparam prom_inst_0.INIT_RAM_3B = 256'h00783030307000CC003C18181838C67C007830303070003800783030307000E0;
defparam prom_inst_0.INIT_RAM_3C = 256'h0078CCCC78001C000078CCCC7800E00000CCCCCCF800F8000078CC7C0CD870D8;
defparam prom_inst_0.INIT_RAM_3D = 256'h001818007E0018180078CCCC7800CC000078CCCC7800DC760078CCCC7800CC78;
defparam prom_inst_0.INIT_RAM_3E = 256'h007ECCCCCC00CC78007ECCCCCC001C00007ECCCCCC00E000603C767E6E3C0600;
defparam prom_inst_0.INIT_RAM_3F = 256'hF80C7CCCCC00CC0000607C667C600000F80C7CCCCC001C00007ECCCCCC00CC00;

endmodule //font8x8
